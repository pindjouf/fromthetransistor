module TxUnit(
    input data_in,


    output data_tx,
    output active,
    output done
    );

endmodule
