module blink (
    input clk,
    output led
);
    
    assign led = clk;
    
endmodule
