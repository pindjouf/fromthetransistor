module design();
    
endmodule
